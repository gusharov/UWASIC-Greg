`default_nettype none



module spi (  
    input clk, sdi, cs,    
    output sdo
);

    
endmodule