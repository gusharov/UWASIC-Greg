`default_nettype none



module spi (  
    input sclk, sdi, cs,    
    output sdo
);

    
endmodule