/*
 * Copyright (c) 2024 Gregory Usharov
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_uwasic_onboarding_Gregory_Usharov (
    
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset

);


    wire [7:0] en_reg_out_7_0;
    wire [7:0] en_reg_out_15_8;
    wire [7:0] en_reg_pwm_7_0;
    wire [7:0] en_reg_pwm_15_8;
    wire [7:0] pwm_duty_cycle;

  pwm_peripheral pwm_peripheral_inst (
      .clk(clk),
      .rst_n(rst_n),
      .en_reg_out_7_0(en_reg_out_7_0),
      .en_reg_out_15_8(en_reg_out_15_8),
      .en_reg_pwm_7_0(en_reg_pwm_7_0),
      .en_reg_pwm_15_8(en_reg_pwm_15_8),
      .pwm_duty_cycle(pwm_duty_cycle),
      .out({uio_out, uo_out})
    );

  wire nuuh;
  spi spi_inst(
    .clk(clk),
    .sclk(ui_in[0]),
    .sdi(ui_in[1]),
    .cs(ui_in[2]),
    .sdo(nuuh),
    .rst_n(rst_n),
    .reg1(en_reg_out_7_0),
    .reg2(en_reg_out_15_8),
    .reg3(en_reg_pwm_7_0),
    .reg4(en_reg_pwm_15_8),
    .reg5(pwm_duty_cycle)
  );
  wire _unused = &{ena, clk, rst_n, ui_in[7:3], uio_in, 1'b0, nuuh};


  // All output pins must be assigned. If not used, assign to 0.
  assign uio_oe = 8'hFF;

  // List all unused inputs to prevent warnings
endmodule
